
`timescale 1ns / 1ps
 
// Design Name: EXAMPLE (13) --->>   Write Verilog code for a 4-bit unsigned up counter with an asynchronous load from the primary input.

module Example13(counter, Input, clk, load);

output [3:0]counter;
input [3:0] Input;
input clk, load;
reg [3:0]counter_reg;

always @(posedge clk or posedge load)
begin
if(load)
counter_reg <= Input;
else 
counter_reg <= counter_reg + 4'b0001;
end

assign counter = counter_reg;

endmodule